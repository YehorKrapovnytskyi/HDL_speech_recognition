package test_package;

    import "DPI-C" function real my_cos(input real x);
    import "DPI-C" function real my_sin(input real x);

    import "DPI-C" function real frand();

endpackage : test_package